module main ( input [1:0] J1, output D5 );

endmodule
