module main ( input [3:0] J1, output D5 );

assign D5 = &J1;

endmodule
